** Generated for: hspiceD
** Generated on: May  1 23:47:05 2022
** Design library name: Analog_test
** Design cell name: TEST_DIFAMP2
** Design view name: schematic
.PARAM cf=200n l1=200n l2=200n l3=200n l4=200n l5=200n  mcap=200n n1=1 n2=1 n3=1  w1=200n w2=200n w3=200n w4=200n w5=200n res=1e3 
+    vstep=1m vocm=0.9 vout=0.9 vdd=1.8 vin=0


.LIB "/home/kmcho/Analog_GPU_RL_SJPark_coop/Eureka_Development/Eureka_Analog_Sizing/eureka/hspice/lib_files/corner_HL18G.lib" ttt

.PROBE TRAN
+    V(op5)
+    V(on4)
+    V(op4)
+    V(on3)
+    V(op3)
+    V(on)
+    V(op)
+    V(op2)
+    V(vdd2)
+    I(v5)
.PROBE AC
+    VDB(on4) VP(on4)
+    VDB(op4) VP(op4)
+    VDB(on3) VP(on3)
+    VDB(op3) VP(op3)
+    VDB(on) VP(on)
+    VDB(op) VP(op)
+    VDB(op2) VP(op2)
.PROBE NOISE
+    V(on4) VP(on4)
+    V(op4) VP(op4)
+    V(on3) VP(on3)
+    V(op3) VP(op3)
+    V(on) VP(on)
+    V(op) VP(op)
+    V(op2) VP(op2)

.NOISE V(op3, on3) v3 1
+    listfreq=1G
.AC DEC 10 10e-3 1e9
.TRAN 10e-9 1e-6 START=0.0

.TEMP 25.0
.OPTION
+    ARTIST=2
+    INGOLD=2
+    PARHIER=LOCAL
+    PSF=2
+    DCON = -1
+    CONV = -1
+    METHOD = GEAR
+    ACCURATE = 1

.param settling_range = 0.1

.measure AC UGF when VDB(op, on) = 0 cross = 1
.measure AC phase_0dB find VP(op, on) when VDB(op, on) = 0
.measure AC PM = param('180+phase_0dB')
.measure AC DC_Gain find VDB(op, on) at=10e-3
.measure AC CM_Gain find VDB(op2) at=10e-3
.measure AC PW_Gain find VDB(op3) at=10e-3
.measure AC CMRR = param('DC_Gain - CM_Gain')
.measure AC PSRR = param('DC_Gain - PW_Gain')

.measure TRAN VH find V(op) at = 2.5e-7
.measure TRAN VL find V(op) at = 7.5e-7 
.measure TRAN OS = param('VH-VL')

.measure TRAN Upper find V(OP5) at = 0
.measure TRAN init find V(OP4) at = 0 
.measure TRAN Upper_bound param('Upper+settling_range*(Upper-init)')
.measure TRAN Lower_bound param('Upper-settling_range*(Upper-init)')

.measure TRAN Upper_trig 
+trig V(OP4) = Upper cross = 1
+targ V(OP4) = Upper_bound cross = last
.measure TRAN Lower_trig
+trig V(OP4) = Lower_bound cross = 1
+targ V(OP4) = Lower_bound cross = last

.measure TRAN I_vdd find I(v5) at = 0
.measure TRAN V_vdd find V(vdd2) at = 0
.measure TRAN pwr = param('(-1)*V_vdd*I_vdd')


** Library name: Analog_180nm
** Cell name: OTA
** View name: schematic
.subckt OTA gnd inn inp outn outp vdd vocm
mpm12 vbp vbp vdd vdd pch_tn w=w4 l=l4 ad='w4<419.5e-9?(int(int(1)/2)*(176.4e-15+w4*200e-9)+(int(1)/2-int(int(1)/2)!=0?176.4e-15+w4*100e-9:0))/1:(int(int(1)/2)*(540e-9*w4)+(int(1)/2-int(int(1)/2)!=0?480e-9*w4:0))/1' as='w4<419.5e-9?(((176.4e-15+w4*100e-9)+int((int(1)-1)/2)*(176.4e-15+w4*200e-9))+(int(1)/2-int(int(1)/2)==0?176.4e-15+w4*100e-9:0))/1:((480e-9*w4+int((int(1)-1)/2)*(540e-9*w4))+(int(1)/2-int(int(1)/2)==0?480e-9*w4:0))/1' pd='w4<419.5e-9?(int(int(1)/2)*2.08e-6+(int(1)/2-int(int(1)/2)!=0?1.88e-6:0))/1:(int(int(1)/2)*(1.08e-6+2*w4)+(int(1)/2-int(int(1)/2)!=0?960e-9+2*w4:0))/1' ps='w4<419.5e-9?((1.88e-6+int((int(1)-1)/2)*2.08e-6)+(int(1)/2-int(int(1)/2)==0?1.88e-6:0))/1:(((960e-9+2*w4)+int((int(1)-1)/2)*(1.08e-6+2*w4))+(int(1)/2-int(int(1)/2)==0?960e-9+2*w4:0))/1' nrd='w4<419.5e-9?(int(int(1)/2)*(176.4e-15+w4*200e-9)+(int(1)/2-int(int(1)/2)!=0?176.4e-15+w4*100e-9:0))/1:((int(int(1)/2)*(540e-9*w4)+(int(1)/2-int(int(1)/2)!=0?480e-9*w4:0))/1)/(w4*w4)'
+nrs='w4<419.5e-9?(((176.4e-15+w4*100e-9)+int((int(1)-1)/2)*(176.4e-15+w4*200e-9))+(int(1)/2-int(int(1)/2)==0?176.4e-15+w4*100e-9:0))/1:(((480e-9*w4+int((int(1)-1)/2)*(540e-9*w4))+(int(1)/2-int(int(1)/2)==0?480e-9*w4:0))/1)/(w4*w4)' m=1
mpm9 net16 vbp vdd vdd pch_tn w=w4 l=l4 ad='w4<419.5e-9?(int(int(1)/2)*(176.4e-15+w4*200e-9)+(int(1)/2-int(int(1)/2)!=0?176.4e-15+w4*100e-9:0))/1:(int(int(1)/2)*(540e-9*w4)+(int(1)/2-int(int(1)/2)!=0?480e-9*w4:0))/1' as='w4<419.5e-9?(((176.4e-15+w4*100e-9)+int((int(1)-1)/2)*(176.4e-15+w4*200e-9))+(int(1)/2-int(int(1)/2)==0?176.4e-15+w4*100e-9:0))/1:((480e-9*w4+int((int(1)-1)/2)*(540e-9*w4))+(int(1)/2-int(int(1)/2)==0?480e-9*w4:0))/1' pd='w4<419.5e-9?(int(int(1)/2)*2.08e-6+(int(1)/2-int(int(1)/2)!=0?1.88e-6:0))/1:(int(int(1)/2)*(1.08e-6+2*w4)+(int(1)/2-int(int(1)/2)!=0?960e-9+2*w4:0))/1' ps='w4<419.5e-9?((1.88e-6+int((int(1)-1)/2)*2.08e-6)+(int(1)/2-int(int(1)/2)==0?1.88e-6:0))/1:(((960e-9+2*w4)+int((int(1)-1)/2)*(1.08e-6+2*w4))+(int(1)/2-int(int(1)/2)==0?960e-9+2*w4:0))/1' nrd='w4<419.5e-9?(int(int(1)/2)*(176.4e-15+w4*200e-9)+(int(1)/2-int(int(1)/2)!=0?176.4e-15+w4*100e-9:0))/1:((int(int(1)/2)*(540e-9*w4)+(int(1)/2-int(int(1)/2)!=0?480e-9*w4:0))/1)/(w4*w4)'
+nrs='w4<419.5e-9?(((176.4e-15+w4*100e-9)+int((int(1)-1)/2)*(176.4e-15+w4*200e-9))+(int(1)/2-int(int(1)/2)==0?176.4e-15+w4*100e-9:0))/1:(((480e-9*w4+int((int(1)-1)/2)*(540e-9*w4))+(int(1)/2-int(int(1)/2)==0?480e-9*w4:0))/1)/(w4*w4)' m='(2*n3)*1'
mpm7 vcmfb net026 net16 net16 pch_tn w=w3 l=l3 ad='w3<419.5e-9?(int(int(1)/2)*(176.4e-15+w3*200e-9)+(int(1)/2-int(int(1)/2)!=0?176.4e-15+w3*100e-9:0))/1:(int(int(1)/2)*(540e-9*w3)+(int(1)/2-int(int(1)/2)!=0?480e-9*w3:0))/1' as='w3<419.5e-9?(((176.4e-15+w3*100e-9)+int((int(1)-1)/2)*(176.4e-15+w3*200e-9))+(int(1)/2-int(int(1)/2)==0?176.4e-15+w3*100e-9:0))/1:((480e-9*w3+int((int(1)-1)/2)*(540e-9*w3))+(int(1)/2-int(int(1)/2)==0?480e-9*w3:0))/1' pd='w3<419.5e-9?(int(int(1)/2)*2.08e-6+(int(1)/2-int(int(1)/2)!=0?1.88e-6:0))/1:(int(int(1)/2)*(1.08e-6+2*w3)+(int(1)/2-int(int(1)/2)!=0?960e-9+2*w3:0))/1' ps='w3<419.5e-9?((1.88e-6+int((int(1)-1)/2)*2.08e-6)+(int(1)/2-int(int(1)/2)==0?1.88e-6:0))/1:(((960e-9+2*w3)+int((int(1)-1)/2)*(1.08e-6+2*w3))+(int(1)/2-int(int(1)/2)==0?960e-9+2*w3:0))/1' nrd='w3<419.5e-9?(int(int(1)/2)*(176.4e-15+w3*200e-9)+(int(1)/2-int(int(1)/2)!=0?176.4e-15+w3*100e-9:0))/1:((int(int(1)/2)*(540e-9*w3)+(int(1)/2-int(int(1)/2)!=0?480e-9*w3:0))/1)/(w3*w3)'
+nrs='w3<419.5e-9?(((176.4e-15+w3*100e-9)+int((int(1)-1)/2)*(176.4e-15+w3*200e-9))+(int(1)/2-int(int(1)/2)==0?176.4e-15+w3*100e-9:0))/1:(((480e-9*w3+int((int(1)-1)/2)*(540e-9*w3))+(int(1)/2-int(int(1)/2)==0?480e-9*w3:0))/1)/(w3*w3)' m='n3*1'
mpm6 net024 vocm net16 net16 pch_tn w=w3 l=l3 ad='w3<419.5e-9?(int(int(1)/2)*(176.4e-15+w3*200e-9)+(int(1)/2-int(int(1)/2)!=0?176.4e-15+w3*100e-9:0))/1:(int(int(1)/2)*(540e-9*w3)+(int(1)/2-int(int(1)/2)!=0?480e-9*w3:0))/1' as='w3<419.5e-9?(((176.4e-15+w3*100e-9)+int((int(1)-1)/2)*(176.4e-15+w3*200e-9))+(int(1)/2-int(int(1)/2)==0?176.4e-15+w3*100e-9:0))/1:((480e-9*w3+int((int(1)-1)/2)*(540e-9*w3))+(int(1)/2-int(int(1)/2)==0?480e-9*w3:0))/1' pd='w3<419.5e-9?(int(int(1)/2)*2.08e-6+(int(1)/2-int(int(1)/2)!=0?1.88e-6:0))/1:(int(int(1)/2)*(1.08e-6+2*w3)+(int(1)/2-int(int(1)/2)!=0?960e-9+2*w3:0))/1' ps='w3<419.5e-9?((1.88e-6+int((int(1)-1)/2)*2.08e-6)+(int(1)/2-int(int(1)/2)==0?1.88e-6:0))/1:(((960e-9+2*w3)+int((int(1)-1)/2)*(1.08e-6+2*w3))+(int(1)/2-int(int(1)/2)==0?960e-9+2*w3:0))/1' nrd='w3<419.5e-9?(int(int(1)/2)*(176.4e-15+w3*200e-9)+(int(1)/2-int(int(1)/2)!=0?176.4e-15+w3*100e-9:0))/1:((int(int(1)/2)*(540e-9*w3)+(int(1)/2-int(int(1)/2)!=0?480e-9*w3:0))/1)/(w3*w3)'
+nrs='w3<419.5e-9?(((176.4e-15+w3*100e-9)+int((int(1)-1)/2)*(176.4e-15+w3*200e-9))+(int(1)/2-int(int(1)/2)==0?176.4e-15+w3*100e-9:0))/1:(((480e-9*w3+int((int(1)-1)/2)*(540e-9*w3))+(int(1)/2-int(int(1)/2)==0?480e-9*w3:0))/1)/(w3*w3)' m='n3*1'
mpm5 outn net13 vdd vdd pch_tn w=w5 l=l5 ad='w5<419.5e-9?(int(int(1)/2)*(176.4e-15+w5*200e-9)+(int(1)/2-int(int(1)/2)!=0?176.4e-15+w5*100e-9:0))/1:(int(int(1)/2)*(540e-9*w5)+(int(1)/2-int(int(1)/2)!=0?480e-9*w5:0))/1' as='w5<419.5e-9?(((176.4e-15+w5*100e-9)+int((int(1)-1)/2)*(176.4e-15+w5*200e-9))+(int(1)/2-int(int(1)/2)==0?176.4e-15+w5*100e-9:0))/1:((480e-9*w5+int((int(1)-1)/2)*(540e-9*w5))+(int(1)/2-int(int(1)/2)==0?480e-9*w5:0))/1' pd='w5<419.5e-9?(int(int(1)/2)*2.08e-6+(int(1)/2-int(int(1)/2)!=0?1.88e-6:0))/1:(int(int(1)/2)*(1.08e-6+2*w5)+(int(1)/2-int(int(1)/2)!=0?960e-9+2*w5:0))/1' ps='w5<419.5e-9?((1.88e-6+int((int(1)-1)/2)*2.08e-6)+(int(1)/2-int(int(1)/2)==0?1.88e-6:0))/1:(((960e-9+2*w5)+int((int(1)-1)/2)*(1.08e-6+2*w5))+(int(1)/2-int(int(1)/2)==0?960e-9+2*w5:0))/1' nrd='w5<419.5e-9?(int(int(1)/2)*(176.4e-15+w5*200e-9)+(int(1)/2-int(int(1)/2)!=0?176.4e-15+w5*100e-9:0))/1:((int(int(1)/2)*(540e-9*w5)+(int(1)/2-int(int(1)/2)!=0?480e-9*w5:0))/1)/(w5*w5)'
+nrs='w5<419.5e-9?(((176.4e-15+w5*100e-9)+int((int(1)-1)/2)*(176.4e-15+w5*200e-9))+(int(1)/2-int(int(1)/2)==0?176.4e-15+w5*100e-9:0))/1:(((480e-9*w5+int((int(1)-1)/2)*(540e-9*w5))+(int(1)/2-int(int(1)/2)==0?480e-9*w5:0))/1)/(w5*w5)' m='n1*1'
mpm4 outp net15 vdd vdd pch_tn w=w5 l=l5 ad='w5<419.5e-9?(int(int(1)/2)*(176.4e-15+w5*200e-9)+(int(1)/2-int(int(1)/2)!=0?176.4e-15+w5*100e-9:0))/1:(int(int(1)/2)*(540e-9*w5)+(int(1)/2-int(int(1)/2)!=0?480e-9*w5:0))/1' as='w5<419.5e-9?(((176.4e-15+w5*100e-9)+int((int(1)-1)/2)*(176.4e-15+w5*200e-9))+(int(1)/2-int(int(1)/2)==0?176.4e-15+w5*100e-9:0))/1:((480e-9*w5+int((int(1)-1)/2)*(540e-9*w5))+(int(1)/2-int(int(1)/2)==0?480e-9*w5:0))/1' pd='w5<419.5e-9?(int(int(1)/2)*2.08e-6+(int(1)/2-int(int(1)/2)!=0?1.88e-6:0))/1:(int(int(1)/2)*(1.08e-6+2*w5)+(int(1)/2-int(int(1)/2)!=0?960e-9+2*w5:0))/1' ps='w5<419.5e-9?((1.88e-6+int((int(1)-1)/2)*2.08e-6)+(int(1)/2-int(int(1)/2)==0?1.88e-6:0))/1:(((960e-9+2*w5)+int((int(1)-1)/2)*(1.08e-6+2*w5))+(int(1)/2-int(int(1)/2)==0?960e-9+2*w5:0))/1' nrd='w5<419.5e-9?(int(int(1)/2)*(176.4e-15+w5*200e-9)+(int(1)/2-int(int(1)/2)!=0?176.4e-15+w5*100e-9:0))/1:((int(int(1)/2)*(540e-9*w5)+(int(1)/2-int(int(1)/2)!=0?480e-9*w5:0))/1)/(w5*w5)'
+nrs='w5<419.5e-9?(((176.4e-15+w5*100e-9)+int((int(1)-1)/2)*(176.4e-15+w5*200e-9))+(int(1)/2-int(int(1)/2)==0?176.4e-15+w5*100e-9:0))/1:(((480e-9*w5+int((int(1)-1)/2)*(540e-9*w5))+(int(1)/2-int(int(1)/2)==0?480e-9*w5:0))/1)/(w5*w5)' m='n1*1'
mpm2 net13 vbp vdd vdd pch_tn w=w4 l=l4 ad='w4<419.5e-9?(int(int(1)/2)*(176.4e-15+w4*200e-9)+(int(1)/2-int(int(1)/2)!=0?176.4e-15+w4*100e-9:0))/1:(int(int(1)/2)*(540e-9*w4)+(int(1)/2-int(int(1)/2)!=0?480e-9*w4:0))/1' as='w4<419.5e-9?(((176.4e-15+w4*100e-9)+int((int(1)-1)/2)*(176.4e-15+w4*200e-9))+(int(1)/2-int(int(1)/2)==0?176.4e-15+w4*100e-9:0))/1:((480e-9*w4+int((int(1)-1)/2)*(540e-9*w4))+(int(1)/2-int(int(1)/2)==0?480e-9*w4:0))/1' pd='w4<419.5e-9?(int(int(1)/2)*2.08e-6+(int(1)/2-int(int(1)/2)!=0?1.88e-6:0))/1:(int(int(1)/2)*(1.08e-6+2*w4)+(int(1)/2-int(int(1)/2)!=0?960e-9+2*w4:0))/1' ps='w4<419.5e-9?((1.88e-6+int((int(1)-1)/2)*2.08e-6)+(int(1)/2-int(int(1)/2)==0?1.88e-6:0))/1:(((960e-9+2*w4)+int((int(1)-1)/2)*(1.08e-6+2*w4))+(int(1)/2-int(int(1)/2)==0?960e-9+2*w4:0))/1' nrd='w4<419.5e-9?(int(int(1)/2)*(176.4e-15+w4*200e-9)+(int(1)/2-int(int(1)/2)!=0?176.4e-15+w4*100e-9:0))/1:((int(int(1)/2)*(540e-9*w4)+(int(1)/2-int(int(1)/2)!=0?480e-9*w4:0))/1)/(w4*w4)'
+nrs='w4<419.5e-9?(((176.4e-15+w4*100e-9)+int((int(1)-1)/2)*(176.4e-15+w4*200e-9))+(int(1)/2-int(int(1)/2)==0?176.4e-15+w4*100e-9:0))/1:(((480e-9*w4+int((int(1)-1)/2)*(540e-9*w4))+(int(1)/2-int(int(1)/2)==0?480e-9*w4:0))/1)/(w4*w4)' m='n2*1'
mpm0 net15 vbp vdd vdd pch_tn w=w4 l=l4 ad='w4<419.5e-9?(int(int(1)/2)*(176.4e-15+w4*200e-9)+(int(1)/2-int(int(1)/2)!=0?176.4e-15+w4*100e-9:0))/1:(int(int(1)/2)*(540e-9*w4)+(int(1)/2-int(int(1)/2)!=0?480e-9*w4:0))/1' as='w4<419.5e-9?(((176.4e-15+w4*100e-9)+int((int(1)-1)/2)*(176.4e-15+w4*200e-9))+(int(1)/2-int(int(1)/2)==0?176.4e-15+w4*100e-9:0))/1:((480e-9*w4+int((int(1)-1)/2)*(540e-9*w4))+(int(1)/2-int(int(1)/2)==0?480e-9*w4:0))/1' pd='w4<419.5e-9?(int(int(1)/2)*2.08e-6+(int(1)/2-int(int(1)/2)!=0?1.88e-6:0))/1:(int(int(1)/2)*(1.08e-6+2*w4)+(int(1)/2-int(int(1)/2)!=0?960e-9+2*w4:0))/1' ps='w4<419.5e-9?((1.88e-6+int((int(1)-1)/2)*2.08e-6)+(int(1)/2-int(int(1)/2)==0?1.88e-6:0))/1:(((960e-9+2*w4)+int((int(1)-1)/2)*(1.08e-6+2*w4))+(int(1)/2-int(int(1)/2)==0?960e-9+2*w4:0))/1' nrd='w4<419.5e-9?(int(int(1)/2)*(176.4e-15+w4*200e-9)+(int(1)/2-int(int(1)/2)!=0?176.4e-15+w4*100e-9:0))/1:((int(int(1)/2)*(540e-9*w4)+(int(1)/2-int(int(1)/2)!=0?480e-9*w4:0))/1)/(w4*w4)'
+nrs='w4<419.5e-9?(((176.4e-15+w4*100e-9)+int((int(1)-1)/2)*(176.4e-15+w4*200e-9))+(int(1)/2-int(int(1)/2)==0?176.4e-15+w4*100e-9:0))/1:(((480e-9*w4+int((int(1)-1)/2)*(540e-9*w4))+(int(1)/2-int(int(1)/2)==0?480e-9*w4:0))/1)/(w4*w4)' m='n2*1'
mnm13 vbp vbn gnd gnd nch_tn w=w1 l=l1 ad='w1<419.5e-9?(int(int(1)/2)*(176.4e-15+w1*200e-9)+(int(1)/2-int(int(1)/2)!=0?176.4e-15+w1*100e-9:0))/1:(int(int(1)/2)*(540e-9*w1)+(int(1)/2-int(int(1)/2)!=0?480e-9*w1:0))/1' as='w1<419.5e-9?(((176.4e-15+w1*100e-9)+int((int(1)-1)/2)*(176.4e-15+w1*200e-9))+(int(1)/2-int(int(1)/2)==0?176.4e-15+w1*100e-9:0))/1:((480e-9*w1+int((int(1)-1)/2)*(540e-9*w1))+(int(1)/2-int(int(1)/2)==0?480e-9*w1:0))/1' pd='w1<419.5e-9?(int(int(1)/2)*2.08e-6+(int(1)/2-int(int(1)/2)!=0?1.88e-6:0))/1:(int(int(1)/2)*(1.08e-6+2*w1)+(int(1)/2-int(int(1)/2)!=0?960e-9+2*w1:0))/1' ps='w1<419.5e-9?((1.88e-6+int((int(1)-1)/2)*2.08e-6)+(int(1)/2-int(int(1)/2)==0?1.88e-6:0))/1:(((960e-9+2*w1)+int((int(1)-1)/2)*(1.08e-6+2*w1))+(int(1)/2-int(int(1)/2)==0?960e-9+2*w1:0))/1' nrd='w1<419.5e-9?(int(int(1)/2)*(176.4e-15+w1*200e-9)+(int(1)/2-int(int(1)/2)!=0?176.4e-15+w1*100e-9:0))/1:((int(int(1)/2)*(540e-9*w1)+(int(1)/2-int(int(1)/2)!=0?480e-9*w1:0))/1)/(w1*w1)'
+nrs='w1<419.5e-9?(((176.4e-15+w1*100e-9)+int((int(1)-1)/2)*(176.4e-15+w1*200e-9))+(int(1)/2-int(int(1)/2)==0?176.4e-15+w1*100e-9:0))/1:(((480e-9*w1+int((int(1)-1)/2)*(540e-9*w1))+(int(1)/2-int(int(1)/2)==0?480e-9*w1:0))/1)/(w1*w1)' m=1
mnm11 vbn vbn gnd gnd nch_tn w=w1 l=l1 ad='w1<419.5e-9?(int(int(1)/2)*(176.4e-15+w1*200e-9)+(int(1)/2-int(int(1)/2)!=0?176.4e-15+w1*100e-9:0))/1:(int(int(1)/2)*(540e-9*w1)+(int(1)/2-int(int(1)/2)!=0?480e-9*w1:0))/1' as='w1<419.5e-9?(((176.4e-15+w1*100e-9)+int((int(1)-1)/2)*(176.4e-15+w1*200e-9))+(int(1)/2-int(int(1)/2)==0?176.4e-15+w1*100e-9:0))/1:((480e-9*w1+int((int(1)-1)/2)*(540e-9*w1))+(int(1)/2-int(int(1)/2)==0?480e-9*w1:0))/1' pd='w1<419.5e-9?(int(int(1)/2)*2.08e-6+(int(1)/2-int(int(1)/2)!=0?1.88e-6:0))/1:(int(int(1)/2)*(1.08e-6+2*w1)+(int(1)/2-int(int(1)/2)!=0?960e-9+2*w1:0))/1' ps='w1<419.5e-9?((1.88e-6+int((int(1)-1)/2)*2.08e-6)+(int(1)/2-int(int(1)/2)==0?1.88e-6:0))/1:(((960e-9+2*w1)+int((int(1)-1)/2)*(1.08e-6+2*w1))+(int(1)/2-int(int(1)/2)==0?960e-9+2*w1:0))/1' nrd='w1<419.5e-9?(int(int(1)/2)*(176.4e-15+w1*200e-9)+(int(1)/2-int(int(1)/2)!=0?176.4e-15+w1*100e-9:0))/1:((int(int(1)/2)*(540e-9*w1)+(int(1)/2-int(int(1)/2)!=0?480e-9*w1:0))/1)/(w1*w1)'
+nrs='w1<419.5e-9?(((176.4e-15+w1*100e-9)+int((int(1)-1)/2)*(176.4e-15+w1*200e-9))+(int(1)/2-int(int(1)/2)==0?176.4e-15+w1*100e-9:0))/1:(((480e-9*w1+int((int(1)-1)/2)*(540e-9*w1))+(int(1)/2-int(int(1)/2)==0?480e-9*w1:0))/1)/(w1*w1)' m=1
mnm10 vcmfb vcmfb gnd gnd nch_tn w=w1 l=l1 ad='w1<419.5e-9?(int(int(1)/2)*(176.4e-15+w1*200e-9)+(int(1)/2-int(int(1)/2)!=0?176.4e-15+w1*100e-9:0))/1:(int(int(1)/2)*(540e-9*w1)+(int(1)/2-int(int(1)/2)!=0?480e-9*w1:0))/1' as='w1<419.5e-9?(((176.4e-15+w1*100e-9)+int((int(1)-1)/2)*(176.4e-15+w1*200e-9))+(int(1)/2-int(int(1)/2)==0?176.4e-15+w1*100e-9:0))/1:((480e-9*w1+int((int(1)-1)/2)*(540e-9*w1))+(int(1)/2-int(int(1)/2)==0?480e-9*w1:0))/1' pd='w1<419.5e-9?(int(int(1)/2)*2.08e-6+(int(1)/2-int(int(1)/2)!=0?1.88e-6:0))/1:(int(int(1)/2)*(1.08e-6+2*w1)+(int(1)/2-int(int(1)/2)!=0?960e-9+2*w1:0))/1' ps='w1<419.5e-9?((1.88e-6+int((int(1)-1)/2)*2.08e-6)+(int(1)/2-int(int(1)/2)==0?1.88e-6:0))/1:(((960e-9+2*w1)+int((int(1)-1)/2)*(1.08e-6+2*w1))+(int(1)/2-int(int(1)/2)==0?960e-9+2*w1:0))/1' nrd='w1<419.5e-9?(int(int(1)/2)*(176.4e-15+w1*200e-9)+(int(1)/2-int(int(1)/2)!=0?176.4e-15+w1*100e-9:0))/1:((int(int(1)/2)*(540e-9*w1)+(int(1)/2-int(int(1)/2)!=0?480e-9*w1:0))/1)/(w1*w1)'
+nrs='w1<419.5e-9?(((176.4e-15+w1*100e-9)+int((int(1)-1)/2)*(176.4e-15+w1*200e-9))+(int(1)/2-int(int(1)/2)==0?176.4e-15+w1*100e-9:0))/1:(((480e-9*w1+int((int(1)-1)/2)*(540e-9*w1))+(int(1)/2-int(int(1)/2)==0?480e-9*w1:0))/1)/(w1*w1)' m='n3*1'
mnm9 net024 net024 gnd gnd nch_tn w=w1 l=l1 ad='w1<419.5e-9?(int(int(1)/2)*(176.4e-15+w1*200e-9)+(int(1)/2-int(int(1)/2)!=0?176.4e-15+w1*100e-9:0))/1:(int(int(1)/2)*(540e-9*w1)+(int(1)/2-int(int(1)/2)!=0?480e-9*w1:0))/1' as='w1<419.5e-9?(((176.4e-15+w1*100e-9)+int((int(1)-1)/2)*(176.4e-15+w1*200e-9))+(int(1)/2-int(int(1)/2)==0?176.4e-15+w1*100e-9:0))/1:((480e-9*w1+int((int(1)-1)/2)*(540e-9*w1))+(int(1)/2-int(int(1)/2)==0?480e-9*w1:0))/1' pd='w1<419.5e-9?(int(int(1)/2)*2.08e-6+(int(1)/2-int(int(1)/2)!=0?1.88e-6:0))/1:(int(int(1)/2)*(1.08e-6+2*w1)+(int(1)/2-int(int(1)/2)!=0?960e-9+2*w1:0))/1' ps='w1<419.5e-9?((1.88e-6+int((int(1)-1)/2)*2.08e-6)+(int(1)/2-int(int(1)/2)==0?1.88e-6:0))/1:(((960e-9+2*w1)+int((int(1)-1)/2)*(1.08e-6+2*w1))+(int(1)/2-int(int(1)/2)==0?960e-9+2*w1:0))/1' nrd='w1<419.5e-9?(int(int(1)/2)*(176.4e-15+w1*200e-9)+(int(1)/2-int(int(1)/2)!=0?176.4e-15+w1*100e-9:0))/1:((int(int(1)/2)*(540e-9*w1)+(int(1)/2-int(int(1)/2)!=0?480e-9*w1:0))/1)/(w1*w1)'
+nrs='w1<419.5e-9?(((176.4e-15+w1*100e-9)+int((int(1)-1)/2)*(176.4e-15+w1*200e-9))+(int(1)/2-int(int(1)/2)==0?176.4e-15+w1*100e-9:0))/1:(((480e-9*w1+int((int(1)-1)/2)*(540e-9*w1))+(int(1)/2-int(int(1)/2)==0?480e-9*w1:0))/1)/(w1*w1)' m='n3*1'
mnm8 outn vbn gnd gnd nch_tn w=w1 l=l1 ad='w1<419.5e-9?(int(int(1)/2)*(176.4e-15+w1*200e-9)+(int(1)/2-int(int(1)/2)!=0?176.4e-15+w1*100e-9:0))/1:(int(int(1)/2)*(540e-9*w1)+(int(1)/2-int(int(1)/2)!=0?480e-9*w1:0))/1' as='w1<419.5e-9?(((176.4e-15+w1*100e-9)+int((int(1)-1)/2)*(176.4e-15+w1*200e-9))+(int(1)/2-int(int(1)/2)==0?176.4e-15+w1*100e-9:0))/1:((480e-9*w1+int((int(1)-1)/2)*(540e-9*w1))+(int(1)/2-int(int(1)/2)==0?480e-9*w1:0))/1' pd='w1<419.5e-9?(int(int(1)/2)*2.08e-6+(int(1)/2-int(int(1)/2)!=0?1.88e-6:0))/1:(int(int(1)/2)*(1.08e-6+2*w1)+(int(1)/2-int(int(1)/2)!=0?960e-9+2*w1:0))/1' ps='w1<419.5e-9?((1.88e-6+int((int(1)-1)/2)*2.08e-6)+(int(1)/2-int(int(1)/2)==0?1.88e-6:0))/1:(((960e-9+2*w1)+int((int(1)-1)/2)*(1.08e-6+2*w1))+(int(1)/2-int(int(1)/2)==0?960e-9+2*w1:0))/1' nrd='w1<419.5e-9?(int(int(1)/2)*(176.4e-15+w1*200e-9)+(int(1)/2-int(int(1)/2)!=0?176.4e-15+w1*100e-9:0))/1:((int(int(1)/2)*(540e-9*w1)+(int(1)/2-int(int(1)/2)!=0?480e-9*w1:0))/1)/(w1*w1)'
+nrs='w1<419.5e-9?(((176.4e-15+w1*100e-9)+int((int(1)-1)/2)*(176.4e-15+w1*200e-9))+(int(1)/2-int(int(1)/2)==0?176.4e-15+w1*100e-9:0))/1:(((480e-9*w1+int((int(1)-1)/2)*(540e-9*w1))+(int(1)/2-int(int(1)/2)==0?480e-9*w1:0))/1)/(w1*w1)' m='n1*1'
mnm7 outp vbn gnd gnd nch_tn w=w1 l=l1 ad='w1<419.5e-9?(int(int(1)/2)*(176.4e-15+w1*200e-9)+(int(1)/2-int(int(1)/2)!=0?176.4e-15+w1*100e-9:0))/1:(int(int(1)/2)*(540e-9*w1)+(int(1)/2-int(int(1)/2)!=0?480e-9*w1:0))/1' as='w1<419.5e-9?(((176.4e-15+w1*100e-9)+int((int(1)-1)/2)*(176.4e-15+w1*200e-9))+(int(1)/2-int(int(1)/2)==0?176.4e-15+w1*100e-9:0))/1:((480e-9*w1+int((int(1)-1)/2)*(540e-9*w1))+(int(1)/2-int(int(1)/2)==0?480e-9*w1:0))/1' pd='w1<419.5e-9?(int(int(1)/2)*2.08e-6+(int(1)/2-int(int(1)/2)!=0?1.88e-6:0))/1:(int(int(1)/2)*(1.08e-6+2*w1)+(int(1)/2-int(int(1)/2)!=0?960e-9+2*w1:0))/1' ps='w1<419.5e-9?((1.88e-6+int((int(1)-1)/2)*2.08e-6)+(int(1)/2-int(int(1)/2)==0?1.88e-6:0))/1:(((960e-9+2*w1)+int((int(1)-1)/2)*(1.08e-6+2*w1))+(int(1)/2-int(int(1)/2)==0?960e-9+2*w1:0))/1' nrd='w1<419.5e-9?(int(int(1)/2)*(176.4e-15+w1*200e-9)+(int(1)/2-int(int(1)/2)!=0?176.4e-15+w1*100e-9:0))/1:((int(int(1)/2)*(540e-9*w1)+(int(1)/2-int(int(1)/2)!=0?480e-9*w1:0))/1)/(w1*w1)'
+nrs='w1<419.5e-9?(((176.4e-15+w1*100e-9)+int((int(1)-1)/2)*(176.4e-15+w1*200e-9))+(int(1)/2-int(int(1)/2)==0?176.4e-15+w1*100e-9:0))/1:(((480e-9*w1+int((int(1)-1)/2)*(540e-9*w1))+(int(1)/2-int(int(1)/2)==0?480e-9*w1:0))/1)/(w1*w1)' m='n1*1'
mnm2 net13 inn net05 gnd nch_tn w=w2 l=l2 ad='w2<419.5e-9?(int(int(1)/2)*(176.4e-15+w2*200e-9)+(int(1)/2-int(int(1)/2)!=0?176.4e-15+w2*100e-9:0))/1:(int(int(1)/2)*(540e-9*w2)+(int(1)/2-int(int(1)/2)!=0?480e-9*w2:0))/1' as='w2<419.5e-9?(((176.4e-15+w2*100e-9)+int((int(1)-1)/2)*(176.4e-15+w2*200e-9))+(int(1)/2-int(int(1)/2)==0?176.4e-15+w2*100e-9:0))/1:((480e-9*w2+int((int(1)-1)/2)*(540e-9*w2))+(int(1)/2-int(int(1)/2)==0?480e-9*w2:0))/1' pd='w2<419.5e-9?(int(int(1)/2)*2.08e-6+(int(1)/2-int(int(1)/2)!=0?1.88e-6:0))/1:(int(int(1)/2)*(1.08e-6+2*w2)+(int(1)/2-int(int(1)/2)!=0?960e-9+2*w2:0))/1' ps='w2<419.5e-9?((1.88e-6+int((int(1)-1)/2)*2.08e-6)+(int(1)/2-int(int(1)/2)==0?1.88e-6:0))/1:(((960e-9+2*w2)+int((int(1)-1)/2)*(1.08e-6+2*w2))+(int(1)/2-int(int(1)/2)==0?960e-9+2*w2:0))/1' nrd='w2<419.5e-9?(int(int(1)/2)*(176.4e-15+w2*200e-9)+(int(1)/2-int(int(1)/2)!=0?176.4e-15+w2*100e-9:0))/1:((int(int(1)/2)*(540e-9*w2)+(int(1)/2-int(int(1)/2)!=0?480e-9*w2:0))/1)/(w2*w2)'
+nrs='w2<419.5e-9?(((176.4e-15+w2*100e-9)+int((int(1)-1)/2)*(176.4e-15+w2*200e-9))+(int(1)/2-int(int(1)/2)==0?176.4e-15+w2*100e-9:0))/1:(((480e-9*w2+int((int(1)-1)/2)*(540e-9*w2))+(int(1)/2-int(int(1)/2)==0?480e-9*w2:0))/1)/(w2*w2)' m='n2*1'
mnm1 net05 vcmfb gnd gnd nch_tn w=w1 l=l1 ad='w1<419.5e-9?(int(int(1)/2)*(176.4e-15+w1*200e-9)+(int(1)/2-int(int(1)/2)!=0?176.4e-15+w1*100e-9:0))/1:(int(int(1)/2)*(540e-9*w1)+(int(1)/2-int(int(1)/2)!=0?480e-9*w1:0))/1' as='w1<419.5e-9?(((176.4e-15+w1*100e-9)+int((int(1)-1)/2)*(176.4e-15+w1*200e-9))+(int(1)/2-int(int(1)/2)==0?176.4e-15+w1*100e-9:0))/1:((480e-9*w1+int((int(1)-1)/2)*(540e-9*w1))+(int(1)/2-int(int(1)/2)==0?480e-9*w1:0))/1' pd='w1<419.5e-9?(int(int(1)/2)*2.08e-6+(int(1)/2-int(int(1)/2)!=0?1.88e-6:0))/1:(int(int(1)/2)*(1.08e-6+2*w1)+(int(1)/2-int(int(1)/2)!=0?960e-9+2*w1:0))/1' ps='w1<419.5e-9?((1.88e-6+int((int(1)-1)/2)*2.08e-6)+(int(1)/2-int(int(1)/2)==0?1.88e-6:0))/1:(((960e-9+2*w1)+int((int(1)-1)/2)*(1.08e-6+2*w1))+(int(1)/2-int(int(1)/2)==0?960e-9+2*w1:0))/1' nrd='w1<419.5e-9?(int(int(1)/2)*(176.4e-15+w1*200e-9)+(int(1)/2-int(int(1)/2)!=0?176.4e-15+w1*100e-9:0))/1:((int(int(1)/2)*(540e-9*w1)+(int(1)/2-int(int(1)/2)!=0?480e-9*w1:0))/1)/(w1*w1)'
+nrs='w1<419.5e-9?(((176.4e-15+w1*100e-9)+int((int(1)-1)/2)*(176.4e-15+w1*200e-9))+(int(1)/2-int(int(1)/2)==0?176.4e-15+w1*100e-9:0))/1:(((480e-9*w1+int((int(1)-1)/2)*(540e-9*w1))+(int(1)/2-int(int(1)/2)==0?480e-9*w1:0))/1)/(w1*w1)' m='(2*n2)*1'
mnm0 net15 inp net05 gnd nch_tn w=w2 l=l2 ad='w2<419.5e-9?(int(int(1)/2)*(176.4e-15+w2*200e-9)+(int(1)/2-int(int(1)/2)!=0?176.4e-15+w2*100e-9:0))/1:(int(int(1)/2)*(540e-9*w2)+(int(1)/2-int(int(1)/2)!=0?480e-9*w2:0))/1' as='w2<419.5e-9?(((176.4e-15+w2*100e-9)+int((int(1)-1)/2)*(176.4e-15+w2*200e-9))+(int(1)/2-int(int(1)/2)==0?176.4e-15+w2*100e-9:0))/1:((480e-9*w2+int((int(1)-1)/2)*(540e-9*w2))+(int(1)/2-int(int(1)/2)==0?480e-9*w2:0))/1' pd='w2<419.5e-9?(int(int(1)/2)*2.08e-6+(int(1)/2-int(int(1)/2)!=0?1.88e-6:0))/1:(int(int(1)/2)*(1.08e-6+2*w2)+(int(1)/2-int(int(1)/2)!=0?960e-9+2*w2:0))/1' ps='w2<419.5e-9?((1.88e-6+int((int(1)-1)/2)*2.08e-6)+(int(1)/2-int(int(1)/2)==0?1.88e-6:0))/1:(((960e-9+2*w2)+int((int(1)-1)/2)*(1.08e-6+2*w2))+(int(1)/2-int(int(1)/2)==0?960e-9+2*w2:0))/1' nrd='w2<419.5e-9?(int(int(1)/2)*(176.4e-15+w2*200e-9)+(int(1)/2-int(int(1)/2)!=0?176.4e-15+w2*100e-9:0))/1:((int(int(1)/2)*(540e-9*w2)+(int(1)/2-int(int(1)/2)!=0?480e-9*w2:0))/1)/(w2*w2)'
+nrs='w2<419.5e-9?(((176.4e-15+w2*100e-9)+int((int(1)-1)/2)*(176.4e-15+w2*200e-9))+(int(1)/2-int(int(1)/2)==0?176.4e-15+w2*100e-9:0))/1:(((480e-9*w2+int((int(1)-1)/2)*(540e-9*w2))+(int(1)/2-int(int(1)/2)==0?480e-9*w2:0))/1)/(w2*w2)' m='n2*1'
r3 net14 net15 res
r2 net13 net037 res
r1 outn net026 1e6
r0 outp net026 1e6
c3 outp gnd cf
c2 outn gnd cf
c1 net037 outn mcap
c0 net14 outp mcap
i0 vdd vbn DC=9e-6
.ends OTA
** End of subcircuit definition.


** Library name: Analog_test
** Cell name: TEST_DIFAMP2
** View name: schematic
xi70 gnd op4 istep on4 op4 vdd vocm OTA
xi68 gnd vcm net016 on3 op3 vdd2 vocm OTA
xi69 gnd op5 net08 on5 op5 vdd vocm OTA
xi67 gnd vcm2 vcm2 on2 op2 vdd vocm OTA
xi66 gnd i1 net011 on op vdd vocm OTA
v14 vcm2 0 DC=550e-3 AC 1
v10 vocm 0 DC=vocm
v12 net011 i2 DC=0 AC 1
v2 vcm 0 DC=550e-3
v1 gnd 0 DC=0
v5 vdd2 0 DC=vdd AC 1
v0 vdd 0 DC=vdd
v7 i2 vcm SIN 0 'vdd/2' 1e6 0
v6 vcm i1 SIN 0 'vdd/2' 1e6 0
c13 op4 0 1e-15
c12 on4 0 1e-15
c11 on5 0 1e-15
c10 op5 0 1e-15
c8 op3 0 1e-15
c9 on3 0 1e-15
c3 on 0 1e-15
c2 op 0 1e-15
c4 on2 0 1e-15
c5 op2 0 1e-15
v8 istep vcm PULSE 0 vstep 0 50e-12 50e-12 500e-3 1
v4 net08 vcm DC=vstep
v3 net016 vcm DC=0 
.END
